interface interf(input wire clk);

	logic reset;
	logic[3:0] I_par;
	logic MSB_in;
	logic LSB_in;
	logic s0;
	logic s1;
	logic[3:0] A_par; 	

endinterface
