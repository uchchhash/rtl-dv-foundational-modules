class transaction;

	logic reset;
	rand logic MSB_in;
	rand logic LSB_in;
	logic s0;
	logic s1;
	rand logic[3:0] I_par;
	logic[3:0] A_par;
	rand logic[3:0] num;
   

endclass
