`include "../tb/agent/cntr_transaction.sv"
`include "../tb/agent/cntr_generator.sv"
`include"../tb/agent/cntr_driver.sv"
`include "../tb/agent/cntr_monitor.sv"
`include "../tb/agent/cntr_coverage.sv"
`include "../tb/agent/cntr_agent.sv"
`include "../tb/environment/cntr_scoreboard.sv"
`include "../tb/environment/cntr_environment.sv"
`include "../tb/test_lib/cntr_base_test.sv"
`include "../tb/tb_top/cntr_tb_top.sv"
`include "../tb/tb_top/cntr_interface.sv"
//`include "../rtl/Binary_counter_Ishraq.svp"
