
`include "../rtl/Universal_Shift_Register_Diptangshu.svp"
`include "../verif/tb_top/shiftReg_interface.sv"
`include "../verif/agent/shiftReg_transaction.sv"
`include "../verif/agent/shiftReg_coverage.sv"
`include "../verif/agent/shiftReg_generator.sv"
`include "../verif/agent/shiftReg_monitor.sv"
`include "../verif/agent/shiftReg_driver.sv"
`include "../verif/agent/shiftReg_agent.sv"
`include "../verif/environment/shiftReg_scoreboard.sv"
`include "../verif/environment/shiftReg_environment.sv" 
`include "../verif/test_lib/shiftReg_base_test.sv"
`include "../verif/tb_top/shiftReg_tb_top.sv"





